`include "uvm_macros.svh"

import uvm_pkg::*;

module tb_test;

initial begin
	`uvm_info("RUN_TEST", "Vivado Script Simulation Test", UVM_NONE);
end
	
endmodule
